`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   16:17:30 10/28/2013
// Design Name:   fft_computer
// Module Name:   /home/bill/workspace/EmbeddedSystemDesign/zynq_project-master/zynq_custom_ip/hw/ise/fft_peripheral/testbench.v
// Project Name:  fft_peripheral
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: fft_computer
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testbench;

	// Inputs
	reg i_clk;
	reg i_rst_n;
	reg i_data_valid;
	
	reg i_data_ready;

	// Outputs
	wire o_data_ready;
	wire o_data_valid;
	wire [31:0] o_data;
	reg[15:0] inReal;
	reg[15:0] inImage;
	wire [31:0] i_data={inImage,inReal};
	wire o_valid_fft;
	wire o_valid_multi;
	wire o_valid_dataCtrl;
	// Instantiate the Unit Under Test (UUT)
	fft_computer uut (
		.i_clk(i_clk), 
		.i_rst_n(i_rst_n), 
		.i_data_valid(i_data_valid), 
		.i_data(i_data), 
		.o_data_ready(o_data_ready), 
		.o_data_valid(o_data_valid), 
		.o_data(o_data), 
		.i_data_ready(i_data_ready),
		.o_valid_fft(o_valid_fft),
		.o_valid_multi(o_valid_multi),
		.o_valid_dataCtrl(o_valid_dataCtrl)
	);

	initial begin
		// Initialize Inputs
		i_clk = 0;
		i_rst_n = 0;
		i_data_valid = 0;
		i_data_ready = 0;
		inReal=0;
		inImage=0;

		// Wait 100 ns for global reset to finish
		#100;
		i_data_ready = 1;
		i_rst_n = 1;
		i_data_valid = 1;
        
		// Add stimulus here
#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;


#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

#2 inReal=128;
#2 inReal=127;
#2 inReal=127;
#2 inReal=126;
#2 inReal=125;
#2 inReal=124;
#2 inReal=122;
#2 inReal=120;
#2 inReal=118;
#2 inReal=115;
#2 inReal=112;
#2 inReal=109;
#2 inReal=106;
#2 inReal=102;
#2 inReal=98;
#2 inReal=94;
#2 inReal=90;
#2 inReal=85;
#2 inReal=81;
#2 inReal=76;
#2 inReal=71;
#2 inReal=65;
#2 inReal=60;
#2 inReal=54;
#2 inReal=48;
#2 inReal=43;
#2 inReal=37;
#2 inReal=31;
#2 inReal=24;
#2 inReal=18;
#2 inReal=12;
#2 inReal=6;
#2 inReal=0;
#2 inReal=-6;
#2 inReal=-12;
#2 inReal=-18;
#2 inReal=-24;
#2 inReal=-31;
#2 inReal=-37;
#2 inReal=-43;
#2 inReal=-48;
#2 inReal=-54;
#2 inReal=-60;
#2 inReal=-65;
#2 inReal=-71;
#2 inReal=-76;
#2 inReal=-81;
#2 inReal=-85;
#2 inReal=-90;
#2 inReal=-94;
#2 inReal=-98;
#2 inReal=-102;
#2 inReal=-106;
#2 inReal=-109;
#2 inReal=-112;
#2 inReal=-115;
#2 inReal=-118;
#2 inReal=-120;
#2 inReal=-122;
#2 inReal=-124;
#2 inReal=-125;
#2 inReal=-126;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-127;
#2 inReal=-126;
#2 inReal=-125;
#2 inReal=-124;
#2 inReal=-122;
#2 inReal=-120;
#2 inReal=-118;
#2 inReal=-115;
#2 inReal=-112;
#2 inReal=-109;
#2 inReal=-106;
#2 inReal=-102;
#2 inReal=-98;
#2 inReal=-94;
#2 inReal=-90;
#2 inReal=-85;
#2 inReal=-81;
#2 inReal=-76;
#2 inReal=-71;
#2 inReal=-65;
#2 inReal=-60;
#2 inReal=-54;
#2 inReal=-48;
#2 inReal=-43;
#2 inReal=-37;
#2 inReal=-31;
#2 inReal=-24;
#2 inReal=-18;
#2 inReal=-12;
#2 inReal=-6;
#2 inReal=0;
#2 inReal=6;
#2 inReal=12;
#2 inReal=18;
#2 inReal=24;
#2 inReal=31;
#2 inReal=37;
#2 inReal=43;
#2 inReal=48;
#2 inReal=54;
#2 inReal=60;
#2 inReal=65;
#2 inReal=71;
#2 inReal=76;
#2 inReal=81;
#2 inReal=85;
#2 inReal=90;
#2 inReal=94;
#2 inReal=98;
#2 inReal=102;
#2 inReal=106;
#2 inReal=109;
#2 inReal=112;
#2 inReal=115;
#2 inReal=118;
#2 inReal=120;
#2 inReal=122;
#2 inReal=124;
#2 inReal=125;
#2 inReal=126;
#2 inReal=127;
#2 inReal=127;

	end
	
	always #1 i_clk=~i_clk;
	
	always@(posedge i_clk)
		$display("%d \t %d",$time,o_data);
	
      
endmodule

